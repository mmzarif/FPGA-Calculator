module conv (input JM1222HM_in1, input JM1222HM_in2, input JM1222HM_in3, input JM1222HM_in4, output JM1222HM_out1, 
output JM1222HM_out2, output JM1222HM_out3, output JM1222HM_out4, output JM1222HM_out5, output JM1222HM_out6, output JM1222HM_out7);

a a1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out1);
b b1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out2);
c c1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out3);
d d1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out4);
e e1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out5);
f f1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out6);
g g1(JM1222HM_in1, JM1222HM_in2, JM1222HM_in3, JM1222HM_in4,JM1222HM_out7);

endmodule


